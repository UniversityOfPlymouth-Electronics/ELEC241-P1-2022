module display_controller (
   output logic [7:0] data,
   output logic rs,
   output logic rw,
   output logic e,
   input logic [7:0] ascii_data,
   input logic write,
   input logic clk);
   

 
always_ff @(posedge clk) begin



end
   
   
endmodule
   
